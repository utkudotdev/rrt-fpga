`ifndef POINT_SV
`define POINT_SV

typedef struct packed {
    logic [31:0] x;
    logic [31:0] y;
} point;

`endif
