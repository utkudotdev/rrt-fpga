typedef struct packed {
    logic [31:0] x;
    logic [31:0] y;
} point;
